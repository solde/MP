--
-- Copyright (c) 2017 XXXX, UPC
-- All rights reserved.
-- 

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

package multis_pkg is

subtype st_arb_peticion is std_logic;
subtype st_arb_concesion is std_logic;

end package multis_pkg;
