--
-- Copyright (c) 2017 XXXX, UPC
-- All rights reserved.
-- 

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

package retardos_bus_pkg is

constant ret_bus: time:= 2 ns;

end package retardos_bus_pkg;
