--
-- Copyright (c) 2017 XXXX, UPC
-- All rights reserved.
-- 

library ieee;		
use ieee.std_logic_1164.all;		
use ieee.numeric_std.all;
use work.param_disenyo_pkg.all;
use work.componentes_pkg.all;
--! @image html camino_2.png 

entity camino_mcd is
   port (reloj, pcero, pe_a, pe_b: std_logic;
	ini_a, ini_b: std_logic;
	a, b: in st_dat;
	s: out st_dat;
	ig, meu: out std_logic);
end camino_mcd;

architecture estruc of camino_mcd is
signal mx_a, mx_b, reg_a, reg_b, mx_cam, t_s: st_dat;
signal t_ig, t_meu, mayor: std_logic;

begin





end estruc;
