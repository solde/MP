--
-- Copyright (c) 2017 XXXX, UPC
-- All rights reserved.
-- 

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.param_disenyo_pkg.all;
use work.controlador_pkg.all;
use work.retardos_controlador_pkg.all;
use work.acciones_pkg.all;
use work.procedimientos_controlador_pkg.all;
--! @image html controlador_iden.png 

entity controlador is
port (reloj, pcero: in std_logic;
		arb_pet: out std_logic;
		arb_conc: in std_logic;
--		trans_bus: out std_logic;
		observacion: in std_logic;
		pet: in tp_contro_e;
		s_estado: in tp_contro_cam_estado;
		s_control: out tp_contro_cam_cntl;
		resp: out tp_contro_s;
		resp_m: in tp_cntl_memoria_e;
		pet_m: out tp_cntl_memoria_s;
		identificador: in natural);
end;
  
architecture compor of controlador is

--type tipoestado is (DES0, DES, DESB, CMPETIQ, INI, ESCINI, LEC, PML, PMEA, PMEF, ESPL, ESPEA, ESPEF, ESB, ESCP, HECHOL, HECHOE,
--						PMEX, ESPX, HECHOX);
signal estado, prxestado: tipoestado;

signal derechos_acceso: std_logic;

signal propia: std_logic;
signal s_esta, expulsion: std_logic;

begin
-- identificacion del emisor de la transaccion
propia <= '1' when resp_m.iden = std_logic_vector(to_unsigned(identificador, resp_m.iden'length)) else '0';

-- determinacion de los derechos de acceso al bloque
derechos_acceso <= '1' when (s_estado.AF and s_estado.EST) = '1' else '0';

-- determinar posible expulsion
s_esta <= '1' when (s_estado.EST) = '1' else '0';
expulsion <= not (s_estado.AF) and s_esta;

-- registro de estado
reg_estado: process (reloj, pcero)
variable v_estado: tipoestado;
begin
	if pcero = '1' then
		v_estado := DES0;
	elsif rising_edge(reloj) then
		v_estado := prxestado;										
	end if;
-- asignacion de la variable a la señal, indicando el retardo
	estado <= v_estado after retardo_estado;
end process;    
   
-- logica de proximo estado

   
-- logica de salida


	
end;
