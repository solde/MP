--
-- Copyright (c) 2017 XXXX, UPC
-- All rights reserved.
-- 

library ieee;
use ieee.std_logic_1164.all;

package retardos_inter_proc_cache_pkg is

constant retAND: time := 2 ns;

end package retardos_inter_proc_cache_pkg;
