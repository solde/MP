--
-- Copyright (c) 2017 XXXX, UPC
-- All rights reserved.
-- 

library IEEE;
use IEEE.std_logic_1164.all;

package estado_pkg is

type tipoestado is (ESP, CALC, CALCNI);

end package estado_pkg;

