--
-- Copyright (c) 2017 XXXX, UPC
-- All rights reserved.
-- 

library ieee;
use ieee.std_logic_1164.all;

package retardos_controlador_pkg is

constant retardo_estado: time := 2 ns;
constant retardo_logica_prx_estado: time := 2 ns;
constant retardo_logica_salida: time := 3 ns;

end package retardos_controlador_pkg;
