--
-- Copyright (c) 2017 XXXX, UPC
-- All rights reserved.
-- 

library ieee;
use ieee.std_logic_1164.all;

package retardos_RegDes_pkg is

constant retREGDES: time := 2 ns;

end package retardos_RegDes_pkg;
