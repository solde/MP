--
-- Copyright (c) 2017 XXXX, UPC
-- All rights reserved.
-- 

library ieee;
use ieee.std_logic_1164.all;

package retardos_otros_pkg is

constant ret_reg_pet: time := 2 ns;
constant ret_mux_pet: time := 2 ns;

constant ret_reg_etiq: time := 2 ns;

end package retardos_otros_pkg;
